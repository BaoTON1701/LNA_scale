** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/ac_hbt_13g2.sch
**.subckt ac_hbt_13g2
Vce net2 GND 5
XQ1 Vc Vb GND GND npn13G2 Nx=1
R1 net2 Vc 40k m=1
Vce1 net1 GND dc 0.8 ac 1m
R2 Vb net1 33k m=1
**** begin user architecture code

*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temp=27
.control
save all
op
print Vc Vb I(Vce)
ac dec 10 10k 100meg
meas ac vnom_at FIND Vc AT=100k
let v3db = vnom_at*0.707
meas ac freq_at when Vc=v3db
write ac_hbt_13g2.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
