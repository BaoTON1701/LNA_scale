** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/mc_hbt_13g2_ac.sch
**.subckt mc_hbt_13g2_ac
Vce net2 GND 5
R1 net2 Vc 40k m=1
Vce1 net1 GND dc 0.8 ac 1m
R2 Vb net1 33k m=1
XQ1 Vc Vb GND GND npn13G2 Nx=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temp=27
.param mc_ok = 1

.control
let mc_runs = 1000
let run = 0
shell rm mc_hbt_3dB.csv
***************** LOOP *********************
dowhile run < mc_runs
reset
set run=$&run
save all
ac dec 10 10k 1000meg
meas ac vnom_at FIND Vc AT=100k
let v3db = vnom_at*0.707
meas ac freq_3dB when Vc=v3db
print freq_3dB >> mc_hbt_3dB.csv
let run=run+1
end
***************** LOOP *********************
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
