** sch_path: /foss/designs/simulations/LNA_design_ihp_test.sch
**.subckt LNA_design_ihp_test
VCC VDD GND 3.3
R2 VDD net2 {Rc} m=1
VCM net1 GND 1.65
E1 net4 net5 VOL=' 'sin(2*3.14*100*time)' '
* noconn #net4
* noconn #net5
V1 net3 net1 0.5 ac 1
XQ1 net2 net3 GND GND npn13G2v Nx=1 El=2.5e-6
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temper = 27
.param vin = 0.05
.param Rc = 875
.temp {temper}
.op
.control
tran 100p 500n
;ac dec 10 10 1Meg

plot vout


.endc


.save all


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
