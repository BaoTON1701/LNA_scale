** sch_path: /foss/designs/simulations/try.sch
**.subckt try
XQ2 net2 net1 GND GND npn13G2l Nx={Nx_var} El={El_var}
V1 VDD GND 3.3
Vib_l VDD net1 0
Vic_l VDD net2 0
xQ1 net4 net3 GND GND npn13G2 Nx={Nx_var}
Vib VDD net3 0
Vic VDD net4 0
Vib_v VDD net5 0
Vic_v VDD net6 0
XQ4 net6 net5 GND GND npn13G2v Nx=1
**** begin user architecture code


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ

.param El_var = 1 temper = 27 Nx_var = 1
.temp {temper}
.op
.control
;control of changing params Nx (number of emitter in a row)
set plotib = ' ';
set plotib_l = ' ';
set plotib_v = ' ';
set plotic = ' ';
set plotic_l = ' ';
set plotic_v = ' ';
set plotbeta = ' ';
set plotbeta_v = ' ';
set plotbeta_l = ' ';
let Nx_1 = 1

repeat 10;
	alterparam Nx_var = $&Nx_1
	reset
	dc V1 0.1 1.6 0.05
	set plotib_l = ( $plotib_l ({$curplot}.I(Vib_l)) );
	set plotic_l = ( $plotic_l ({$curplot}.I(Vic_l)) );
	set plotbeta_l = ( $plotbeta_l {$curplot}.I(vic_l)/{$curplot}.I(vib_l) );
	set plotib_v = ( $plotib_v ({$curplot}.I(Vib_v)) );
	set plotic_v = ( $plotic_v ({$curplot}.I(Vic_v)) );
	set plotbeta_v = ( $plotbeta_v {$curplot}.I(vic_v)/{$curplot}.I(vib_v) );
	set plotib =   ( $plotib ({$curplot}.I(Vib)) );
	set plotic =   ( $plotic   ({$curplot}.I(Vic)) );
	set plotbeta =   ( $plotbeta {$curplot}.I(vic)/{$curplot}.I(vib) );
	let Nx_1 = Nx_1 + 1
end;

plot loglog $plotib $plotib_l $plotib_v;
plot loglog $plotic $plotic_l $plotic_v;
plot loglog $plotbeta $plotbeta_l $plotbeta_v;
plot loglog ($plotbeta) vs ($plotic);
;set wr_singlescale;
;set wr_vecnames;
;wrdata gummel_npn13g2_Nx.txt $plotib $plotic $plotbeta;
;wrdata gummel_npn13g2l_Nx.txt $plotib_l $plotic_l $plotbeta_l;
;wrdata gummel_npn13g2v_Nx.txt $plotib_v $plotic_v $plotbeta_v;

.endc

.save all


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
