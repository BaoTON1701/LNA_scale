** sch_path: /foss/designs/simu_test/npn_scaling.sch
**.subckt npn_scaling
XQ2 net10 net1 GND GND npn13G2l Nx={Nx_var} El=1.7
V1 VDD GND 3.3
Vib_l VDD net1 0
Vic_l VDD net10 0
xQ1 net3 net2 GND GND npn13G2 Nx=9
Vib VDD net2 0
Vic VDD net3 0
Vib_v VDD net4 0
Vic_v VDD net5 0
XQ3 net5 net4 GND GND npn13G2v Nx={Nx_var} El={El_var}
* noconn #net9
xQ10 net8 net6 GND GND npn13G2 Nx=10
xQ11 net8 net6 GND GND npn13G2 Nx=10
xQ12 net8 net6 GND GND npn13G2 Nx=10
xQ13 net8 net6 GND GND npn13G2 Nx=10
xQ14 net8 net6 GND GND npn13G2 Nx=7
XQ15 net9 net7 GND GND npn13G2l Nx=4 El=4
XQ16 net9 net7 GND GND npn13G2l Nx=4 El=4
XQ17 net9 net7 GND GND npn13G2l Nx=4 El=4
* noconn #net6
* noconn #net8
* noconn #net7
xQ4 net3 net2 GND GND npn13G2 Nx=9
XQ5 net14 net11 GND GND npn13G2l Nx={Nx_var} El={El_var}
Vib_l1 VDD net11 0
Vic_l1 VDD net14 0
Vib1 VDD net15 0
Vic1 VDD net16 0
Vib_v1 VDD net12 0
Vic_v1 VDD net13 0
XQ7 net13 net12 GND GND npn13G2v Nx={Nx_var} El={El_var}
xQ6 net16 net15 GND GND npn13G2 Nx={Nx_var}
**** begin user architecture code


*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
;Note: Nx of npn13g2 Nx = 1-10
;Nx of npn13g2l Nx = 1-4
;Nx of npn13g2v Nx = 1-8






.param El_var = 1 temper = 27 Nx_var = 1
.param mc_ok = 1
.temp {temper}
.op
.control
echo -----------------------------------------------------
echo starting DC sim
echo -----------------------------------------------------
control of changing params Nx (number of emitter in a row)
set plotib = ' ';
set plotib_l = ' ';
set plotib_v = ' ';
set plotic = ' ';
set plotic_l = ' ';
set plotic_v = ' ';
set plotbeta = ' ';
set plotbeta_v = ' ';
set plotbeta_l = ' ';

set plotib_l1 = ' ';
set plotib_v1 = ' ';
set plotic_l1 = ' ';
set plotic_v1 = ' ';
set plotbeta_v1 = ' ';
set plotbeta_l1 = ' ';

let Nx_1 = 1

repeat 10;
	echo ---------------------------------
	alterparam Nx_var = $&Nx_1
	reset
	op
	dc V1 0.1 1.6 0.05
	if Nx_1 < 5
		set plotib_l = ( $plotib_l ({$curplot}.I(Vib_l1)) );
		set plotic_l = ( $plotic_l ({$curplot}.I(Vic_l1)) );
		set plotbeta_l = ( $plotbeta_l {$curplot}.I(vic_l1)/{$curplot}.I(vib_l1) );
	end;
	if Nx_1 < 9
		set plotib_v = ( $plotib_v ({$curplot}.I(Vib_v1)) );
		set plotic_v = ( $plotic_v ({$curplot}.I(Vic_v1)) );
		set plotbeta_v = ( $plotbeta_v {$curplot}.I(vic_v1)/{$curplot}.I(vib_v1) );
	end;
	set plotib =   ( $plotib ({$curplot}.I(Vib1)) );
	set plotic =   ( $plotic   ({$curplot}.I(Vic1)) );
	set plotbeta =   ( $plotbeta {$curplot}.I(vic1)/{$curplot}.I(vib1) );
	let Nx_1 = Nx_1 + 1
	echo -----------------------------------
end;

let El_1 = 1
repeat 8;
	echo ----------------------------------
	alterparam Nx_Var = 1
	alterparam El_var = $&El_1
	reset
	dc V1 0.1 1.6 0.05
	if El_1 < 2.6
		set plotib_l = ( $plotib_l1 ({$curplot}.I(Vib_l1)) );
		set plotic_l = ( $plotic_l1 ({$curplot}.I(Vic_l1)) );
		set plotbeta_l = ( $plotbeta_l1 {$curplot}.I(vic_l1)/{$curplot}.I(vib_l1) );
	end;
	if El_1 < 5.1
		set plotib_v = ( $plotib_v1 ({$curplot}.I(Vib_v1)) );
		set plotic_v = ( $plotic_v1 ({$curplot}.I(Vic_v1)) );
		set plotbeta_v = ( $plotbeta_v1 {$curplot}.I(vic_v1)/{$curplot}.I(vib_v1) );
	end;
	let El_1 = El_1 + 1
	echo -----------------------------------

set wr_singlescale;
set wr_vecnames;
wrdata gummel_npn13g2_Nx.txt $plotib $plotic $plotbeta;
wrdata gummel_npn13g2l_Nx.txt $plotib_l $plotic_l $plotbeta_l;
wrdata gummel_npn13g2v_Nx.txt $plotib_v $plotic_v $plotbeta_v;

wrdata gummel_npn13g2l_El.txt $plotib_l1 $plotic_l1 $plotbeta_l1;
wrdata gummel_npn13g2v_El.txt $plotib_v1 $plotic_v1 $plotbeta_v1;

.endc


.save all

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
