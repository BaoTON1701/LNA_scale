** sch_path: /foss/designs/simu_test/rlc.sch
**.subckt rlc
R1 A 0 1k m=1
C1 A B 50nF m=1
L1 B C 10mH m=1
E1 C 0 VOL=' '3*cos(time*time*1e6)' '
**** begin user architecture code


.control
tran 10n 10m
;plot v(A) v(C)
.endc
.save all


**** end user architecture code
**.ends
.end
