** sch_path: /foss/designs/simulations/LNA_new.sch
**.subckt LNA_new
V1 VDD GND 2.4
XQ1 net3 vin1 net1 GND npn13G2v Nx=8 El=2.5e-6
XQ2 vout2 vin2 net1 GND npn13G2v Nx=8 El=2.5e-6
I0 net1 GND 4m
R1 VDD vout1 600 m=1
R2 VDD vout2 600 m=1
V2 net2 GND 1.2
E1 vin1 net2 VOL=' '0.005*sin(2*3.14*100000*time)' '
E2 vin2 net2 VOL=' '-0.005*sin(2*pi*100000*time)' '
V3 vout1 net3 0
**** begin user architecture code


.control
tran 1n 100u

plot i(V3)
plot (vin1 - vin2)
.endc
.op
;print @q.xq1.qnpn13g2v[ic] @q.xq1.qnpn13g2v[vce] @q.xq1.qnpn13g2v[vbe]
;print @q.xq2.qnpn13g2v[ic] @q.xq2.qnpn13g2v[vce] @q.xq2.qnpn13g2v[vbe]

.save all



.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
