** sch_path: /foss/designs/simulations/simple_CE_amp.sch
**.subckt simple_CE_amp
XQ1 net1 net2 GND GND npn13G2l Nx=1 El=2.5
V1 net2 in 0.8
E1 in GND VOL=' 0.05*sin(2*3.14*1e5*time) '
R1 VDD out 1k m=1
V2 VDD GND 3.3
VIC out net1 0
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ


.control
	tran 10u 20u
	set nolegend;
	plot (out ) title 'Voltage Gain'
	;plot I(VIC) title 'Ic v. time' ylabel 'Ic'
 	;plot (-I(E1)) title 'Ib v. time' ylabel 'Ib'
	;plot I(VIC)/(-I(E1)) title 'beta v. time'
	;plot I(VIC)/ (in) title 'gm v. time'

.endc
.save all

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
