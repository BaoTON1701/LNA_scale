** sch_path: /foss/designs/simu_test/noise_bipolar.sch
**.subckt noise_bipolar
V1 VDD GND dc 1 ac 1
XQ2 net2 net1 GND GND npn13G2v Nx=4 El=5e-6
VBE net1 GND 0.6
V2 VDD net2 0
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.control
set plot1 = ' ';
let VBE1  = 0.65
repeat 1;
	alter VBE $&VBE1
	noise i(V2) 0 dec 10 1 10MEG
	setplot noise1
	set sqrnoise;
	plot onoise_spectrum
	;set plot1 ( $plot1 {$curplot}.inoise_spectrum );
	let VBE1 = VBE1 + 0.5
end;
.endc
.save all


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
