** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/mc_hbt_13g2.sch
**.subckt mc_hbt_13g2
Vce net3 GND 1.5
I0 GND net1 1u
Vc net3 net2 0
.save i(vc)
XQ1 net2 net1 GND GND npn13G2 Nx=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ_stat
*.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temp=27
.param mc_ok = 1

.control
save all
let mc_runs = 1000
let run = 0
set curplot=new
set scratch=$curplot
setplot $scratch
let Ic=unitvec(mc_runs)

***************** LOOP *********************
dowhile run < mc_runs

op
set run=$&run
set dt=$curplot
setplot $scratch
let out{$run}={$dt}.I(Vc)
let Ic[run]= {$dt}.I(Vc)
setplot $dt
reset
let run=run+1
end
***************** LOOP *********************

wrdata mc_hbt_op.csv {$scratch}.Ic
write mc_hbt_op.raw
echo
print {$scratch}.Ic

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
