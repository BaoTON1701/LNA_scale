** sch_path: /foss/designs/untitled-1.sch
**.subckt untitled-1
XQ1 net1 net2 GND GND npn13G2l Nx=1 El=2.5
V1 net1 GND 0
VBE net2 GND {VBE1}
**** begin user architecture code


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ

.control
	param VBE1=0.4;0.5;0.6
	dc V1 0 1 0.05
	plot all -i(V1)

.endc

.save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
