** sch_path: /foss/designs/simu_test/ihp_bipolar.sch
**.subckt ihp_bipolar
V1 vc GND 0
VBE net1 GND 0.6
XQ2 vc net1 GND GND npn13G2v Nx=1
XQ3 net2 net3 net4 net5 npn13G2l Nx=1 El=2.5
**** begin user architecture code


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temper = -196
.temp {temper};

.control
set plotic = ' ';
set plotib = ' ';
set plotbeta = ' ';

let VBEE = 0.6;

;repeat 5;
;    alter VBE $&VBEE;
;    dc V1 0 1 0.05;
;    set plotic = ( $plotic (-{$curplot}.I(V1)) );
;    set plotib = ( $plotib (-{$curplot}.I(VBE)) );
;    set plotbeta = ( $plotbeta {$curplot}.I(V1)/{$curplot}.I(VBE) );
;    let VBEE = VBEE + 0.05;


;path using array of value instead of step

foreach val1 -196 27
	alterparam temper = $val1
	reset
	let V1 = 3
	dc VBE 0.1 2 0.05
	set plotic = ( $plotic ({$curplot}.I(V1)) );
        set plotib = ( $plotib (-{$curplot}.I(VBE)) );
        set plotbeta = ( $plotbeta {$curplot}.I(V1)/{$curplot}.I(VBE) );
end;

;set nolegend;
set xbrushwidth=2;
plot  $plotic title 'Ic vs VCE' xlabel 'VCE (V)' ylabel 'I_c';
plot  $plotib title 'Ib vs VCE' xlabel 'VCE (V)' ylabel 'I_b';
plot  $plotbeta title 'beta vs VCE' xlabel 'VCE (V)' ylabel 'beta';



.endc
.save all

**** end user architecture code
**.ends
.GLOBAL GND
.end
