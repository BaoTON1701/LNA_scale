** sch_path: /foss/designs/simulations/LNA_design_ihp.sch
**.subckt LNA_design_ihp VCM Vin1 Vin2 Vin1 Vin2 Vout1 Vout2 IEE Vout1 Vout2 VCM IEE
*.opin VCM
*.opin Vin1
*.opin Vin2
*.ipin Vin1
*.ipin Vin2
*.opin Vout1
*.opin Vout2
*.iopin IEE
*.ipin Vout1
*.ipin Vout2
*.ipin VCM
*.opin IEE
VCC VDD GND 3.3
XQ1 Vout1 Vin1 IEE GND npn13G2l Nx=1 El=2.5
R2 VDD Vout1 {Rc} m=1
XQ2 Vout2 Vin2 IEE GND npn13G2l Nx=1 El=2.5
R4 VDD Vout2 {Rc} m=1
VCM VCM GND 1.65
IEE IEE GND 4m
R1 Vout1 GND 1k m=1
R3 Vout2 GND 1k m=1
E1 net3 net4 VOL=' 'sin(2*3.14*100*time)' '
* noconn #net3
* noconn #net4
V1 Vin1 VCM 0.5 ac 1
V2 Vin2 VCM 0.5 ac 1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ



.param temper = 27
.param vin = 0.05
.param Rc = 875
.temp {temper}
.op
.control
tran 100p 500n
;ac dec 10 10 1Meg

plot vout


.endc


.save all


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
