** sch_path: /foss/designs/untitled-5.sch
**.subckt untitled-5
V1 VDD GND 3.3
XQ1 vout1 net4 net1 GND npn13G2v Nx=1 El=2.5e-6
XQ2 vout2 net3 net1 GND npn13G2v Nx=1 El=2.5e-6
I0 net1 GND 4m
R1 VDD vout1 825 m=1
R2 VDD vout2 825 m=1
V2 net2 GND 1.65
E1 net4 net2 VOL=' '0.5*sin(2*3.14*100000*time)' '
E2 net2 net3 VOL=' '0.5*sin(2*pi*100000*time)' '
**** begin user architecture code


.control
tran 1n 10u
plot vout1 vout2
plot vout1 - vout2
.endc
.save all



.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
